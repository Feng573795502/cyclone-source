`timescale 1ns/1ns
module lvds_ip_auto_align_test();


endmodule  